`timescale 1ns / 1ps

package packet_pkg;

 `include "packet_data.sv"
    
endpackage